`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:39:02 11/24/2018
// Design Name:   mips
// Module Name:   C:/Users/Eadral/ISE/P5/mips_tb.v
// Project Name:  P5
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mips
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module mips_tb;

	// Inputs
	reg clk;
	reg reset;

	// Instantiate the Unit Under Test (UUT)
	mips uut (
		.clk(clk), 
		.reset(reset)
	);
	integer i;
	
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;

		// Wait 100 ns for global reset to finish
		#5 clk = ~clk;
		#5 clk = ~clk;
		#5 clk = ~clk;
		reset = 0;
		#5 clk = ~clk;
		
	
		for (i = 0; i < 200; i = i + 1)
			#5 clk = ~clk;
        
		$finish;
	end
      
endmodule

